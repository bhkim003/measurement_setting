//////////////////////////////////////////////////////////////////////////////////
// Engineer: Kim Beomseokfp
// Contact: kimbss470@snu.ac.kr
// 
// Create Date: 16/07/2024 
// Design Name: OpalKelly frontpanel for USB3 in Verilog
// Module Name: DDR3Interface (v2) : do not care single_rate
// Project Name: 2024TapeOut
// Target Devices: XEM7360-K160T
// Tool versions: 2024.1
// Description: Muxing/Demuxing axi signals from/to CHIP/okfp(okFrontPanel) and 
//              connecting to MIG
//
//////////////////////////////////////////////////////////////////////////////////

module DDR3Interface (
    input  wire          sys_clk_p,
    input  wire          sys_clk_n,
    
    input  wire          okRstn,
    input  wire          clk_wiz_locked,

    output wire          clk,         // gen by MIG
    output wire          mig_rstn,    // AND of mig_rstn and clk_wiz_locked
    input  wire          mig_abort,

    inout  wire [ 31:0]  ddr3_dq,
    inout  wire [  3:0]  ddr3_dqs_p,
    inout  wire [  3:0]  ddr3_dqs_n,
    output wire [ 15:0]  ddr3_addr,
    output wire [  2:0]  ddr3_ba,
    output wire          ddr3_ras_n,
    output wire          ddr3_cas_n,
    output wire          ddr3_we_n,
    output wire          ddr3_reset_n,  
    output wire          ddr3_ck_p,
    output wire          ddr3_ck_n,
    output wire          ddr3_cke,
    output wire          ddr3_cs_n,
    output wire          ddr3_odt,
    output wire [  3:0]  ddr3_dm,
    output wire          init_calib_complete,

    input  wire          axi_master, 
    input  wire          chip_store_byte4,    // only write 4byte in the 1st tranfer of the burst
    input  wire          chip_single_rate,
    input  wire [ 27:0]  chip_axi_awaddr,     // Write address
    input  wire [  7:0]  chip_axi_awlen,
    input  wire          chip_axi_awvalid,
    output wire          chip_axi_awready,

    input  wire [255:0]  chip_axi_wdata,      // Write data 
    input  wire          chip_axi_wvalid,
    output wire          chip_axi_wready,

    input  wire [ 27:0]  chip_axi_araddr,     // Read address
    input  wire [  7:0]  chip_axi_arlen,
    input  wire          chip_axi_arvalid,
    output wire          chip_axi_arready,

    output wire [255:0]  chip_axi_rdata,      // Read data
    output wire          chip_axi_rvalid,     // toggled when chip_single_rate == 1'b1
    output wire          chip_axi_rvalid_tmp,
    input  wire          chip_axi_rready,

    input  wire [ 27:0]  okfp_axi_awaddr,     // Write address
    input  wire [  7:0]  okfp_axi_awlen,
    input  wire          okfp_axi_awvalid,
    output wire          okfp_axi_awready,

    input  wire [255:0]  okfp_axi_wdata,      // Write data 
    input  wire          okfp_axi_wvalid,
    output wire          okfp_axi_wready,

    input  wire [ 27:0]  okfp_axi_araddr,     // Read address
    input  wire [  7:0]  okfp_axi_arlen,
    input  wire          okfp_axi_arvalid,
    output wire          okfp_axi_arready,

    output wire [255:0]  okfp_axi_rdata,      // Read data
    output wire          okfp_axi_rvalid,
    input  wire          okfp_axi_rready,

    /* Debug */
    output wire          wstate_debug,
    output wire          s_axi_wready_debug,
    output wire          rstate_debug,
    output wire          s_axi_rready_debug,
    output reg  [ 31:0]  mig_rstate_cnt,
    output reg  [ 31:0]  mig_rvalid_cnt,
    output reg  [ 31:0]  mig_wstate_cnt,
    output reg  [ 31:0]  mig_wvalid_cnt
);

    /* States */
    localparam IDLE  = 2'd0;
    localparam WRITE = 2'd1;
    localparam READ  = 2'd2;


    /* AXI master */
    localparam OKFP = 1'b0;
    localparam CHIP = 1'b1;


    //************************************************************
    //  Wires & Regs
    //************************************************************

    /* AXI interface for MIG */
    wire [27:0]   s_axi_awaddr;
    wire [7:0]    s_axi_awlen;
    wire          s_axi_awvalid;
    wire          s_axi_awready;

    wire [255:0]  s_axi_wdata;
    wire          s_axi_wvalid;
    wire          s_axi_wready;
    reg  [31:0]   s_axi_wstrb;      // generated by DDR3Interface, comb.
    wire          s_axi_wlast;      // generated by DDR3Interface 

    wire          s_axi_bid;
    wire [1:0]    s_axi_bresp;
    wire          s_axi_bvalid;

    wire [27:0]   s_axi_araddr;
    wire [7:0]    s_axi_arlen;
    wire          s_axi_arvalid;
    wire          s_axi_arready;

    wire [255:0]  s_axi_rdata;
    // wire [255:0]  s_axi_rdata_tmp;  // to support single-rate
    // reg  [255:0]  s_axi_rdata_tmp_buf;  // to support single-rate
    wire          s_axi_rlast;
    wire          s_axi_rvalid;
    wire          s_axi_rready;
    wire [1:0]    s_axi_rresp;
    wire          s_axi_rid;


    /* MIG */
    wire rst;
    wire rstn;   
    reg  aresetn;
    wire mmcm_locked;


    /* AXI control */
    reg [1:0]  state;
    wire       wstart;
    wire       rstart;
    wire       wdone;
    wire       rdone;

    reg [31:0] awaddr_buf;
    reg [ 7:0] awlen_buf;
    reg [ 7:0] wcnt;         // write transfer counter

    reg [31:0] araddr_buf;
    reg [ 7:0] arlen_buf;
    reg [ 7:0] rcnt;         // read transfer counter


    /* Self-wstrb-generation */
    reg        chip_store_byte4_buf;


    //************************************************************
    // Generate Reset
    //************************************************************
    assign mig_rstn = ~rst;
    assign rstn = mig_rstn & clk_wiz_locked;


    //************************************************************
    // AXI Crossbar
    //************************************************************
    assign s_axi_awaddr     = (axi_master==CHIP) ? chip_axi_awaddr  : okfp_axi_awaddr;
    assign s_axi_awlen      = (axi_master==CHIP) ? chip_axi_awlen   : okfp_axi_awlen;
    assign s_axi_awvalid    = (axi_master==CHIP) ? chip_axi_awvalid : okfp_axi_awvalid;
    // assign chip_axi_awready = (axi_master==CHIP) ? s_axi_awready : 1'b0;
    // assign okfp_axi_awready = (axi_master==OKFP) ? s_axi_awready : 1'b0; 
    assign chip_axi_awready = (axi_master==CHIP) ? s_axi_awready && (state==IDLE) : 1'b0;
    assign okfp_axi_awready = (axi_master==OKFP) ? s_axi_awready && (state==IDLE) : 1'b0; 

    assign s_axi_wdata      = (axi_master==CHIP) ? chip_axi_wdata  : okfp_axi_wdata;
    assign s_axi_wvalid     = (axi_master==CHIP) ? chip_axi_wvalid : okfp_axi_wvalid;

    // assign chip_axi_wready  = (axi_master==CHIP) ? s_axi_wready : 1'b0;
    // assign okfp_axi_wready  = (axi_master==OKFP) ? s_axi_wready : 1'b0;
    assign chip_axi_wready  = (axi_master==CHIP) ? s_axi_wready & (wstart || (state==WRITE)) : 1'b0;     // wready is valid only when awready is valid, prevent handshaking of wdata from being followed by of awaddr
    assign okfp_axi_wready  = (axi_master==OKFP) ? s_axi_wready & (wstart || (state==WRITE)) : 1'b0;

    assign s_axi_araddr     = (axi_master==CHIP) ? chip_axi_araddr  : okfp_axi_araddr;
    assign s_axi_arlen      = (axi_master==CHIP) ? chip_axi_arlen   : okfp_axi_arlen;
    assign s_axi_arvalid    = (axi_master==CHIP) ? chip_axi_arvalid : okfp_axi_arvalid;
    // assign chip_axi_arready = (axi_master==CHIP) ? s_axi_arready: 1'b0;
    // assign okfp_axi_arready = (axi_master==OKFP) ? s_axi_arready: 1'b0;
    assign chip_axi_arready = (axi_master==CHIP) ? s_axi_arready && (state==IDLE) : 1'b0;
    assign okfp_axi_arready = (axi_master==OKFP) ? s_axi_arready && (state==IDLE) : 1'b0;

    assign chip_axi_rdata   = (axi_master==CHIP) ? s_axi_rdata : 'd0;
    assign okfp_axi_rdata   = (axi_master==OKFP) ? s_axi_rdata : 'd0;
    assign s_axi_rready     = (axi_master==CHIP) ? chip_axi_rready : okfp_axi_rready;
    assign chip_axi_rvalid  = (axi_master==CHIP) ? s_axi_rvalid : 1'b0;
    assign okfp_axi_rvalid  = (axi_master==OKFP) ?  s_axi_rvalid : 1'b0;

    /* Debug */
    assign wstate_debug = wstart || (state==WRITE);
    assign s_axi_wready_debug = s_axi_wready;
    assign rstate_debug = rstart || (state==READ);
    assign s_axi_rready_debug = s_axi_rready;


    //************************************************************
    // Transfer counter 
    //************************************************************
    assign wstart = s_axi_awready & s_axi_awvalid;
    assign rstart = s_axi_arready & s_axi_arvalid;
    assign s_axi_wlast = s_axi_wready && s_axi_wvalid && ((wstart && (s_axi_awlen == 8'd0)) || ((state==WRITE) && (awlen_buf == wcnt))) ;
    assign wdone = (state==WRITE) && s_axi_wlast;
    assign rdone = (state==READ) && s_axi_rlast && s_axi_rready && s_axi_rvalid;


    always @(posedge clk or negedge rstn) begin
        if (~rstn) begin
            state <= IDLE;
        end
        else begin  
            case (state) 
                IDLE: begin
                    if      (rstart) state <= READ;
                    else if (wstart && (!s_axi_wlast)) state <= WRITE;
                    else             state <= IDLE;
                end
                WRITE: begin
                    if (wdone || mig_abort) state <= IDLE;
                    else                    state <= WRITE;
                end
                READ: begin
                    if (rdone || mig_abort) state <= IDLE;
                    else                    state <= READ;
                end
            endcase
        end
    end

    always @(posedge clk or negedge rstn) begin
        if (~rstn) begin
            awaddr_buf <= 32'd0;
            awlen_buf  <= 8'd0;
            wcnt       <= 8'd0;

            araddr_buf <= 32'd0;
            arlen_buf  <= 8'd0;
            rcnt       <= 8'd0;

            mig_rstate_cnt <= 32'd0;
            mig_rvalid_cnt <= 32'd0;
            mig_wstate_cnt <= 32'd0;
            mig_wvalid_cnt <= 32'd0;
        end
        else begin  
            case (state) 
                IDLE: begin
                    // capture addr & len
                    if (wstart) begin
                        awaddr_buf <= s_axi_awaddr;
                        awlen_buf  <= s_axi_awlen;
                        araddr_buf <= 'd0;
                        arlen_buf  <= 'd0;

                        if (axi_master==CHIP) mig_wstate_cnt <= mig_wstate_cnt + 16'd1;
                    end
                    else if (rstart) begin
                        awaddr_buf <= 'd0;
                        awlen_buf  <= 'd0;
                        araddr_buf <= s_axi_araddr;
                        arlen_buf  <= s_axi_arlen;

                        if (axi_master==CHIP) mig_rstate_cnt <= mig_rstate_cnt + 16'd1;
                    end
                    else begin
                        awaddr_buf <= 'd0;
                        awlen_buf  <= 'd0;
                        araddr_buf <= 'd0;
                        arlen_buf  <= 'd0;
                    end

                    // reset wcnt & rcnt
                    if (wstart && s_axi_wready && s_axi_wvalid) begin    // handshake of address and data can be completed simultaneously in AXI-write
                        if (s_axi_wlast) wcnt <= 8'd0;
                        else       wcnt <= wcnt + 8'd1;
                        // wcnt <= wcnt + 8'd1;
                        rcnt <= 8'd0;
                        if (axi_master==CHIP) mig_wvalid_cnt <= mig_wvalid_cnt + 32'd1;
                    end
                    else begin
                        wcnt <= 8'd0;
                        rcnt <= 8'd0;
                    end
                end

                WRITE: begin
                    if (s_axi_wready && s_axi_wvalid) begin
                        if (wdone) wcnt <= 8'd0;
                        else       wcnt <= wcnt + 8'd1;
                        
                        if (axi_master==CHIP) mig_wvalid_cnt <= mig_wvalid_cnt + 32'd1;
                    end

                end

                READ: begin
                    if (s_axi_rready && s_axi_rvalid) begin
                        if (rdone) rcnt <= 8'd0;
                        else       rcnt <= rcnt + 8'd1;

                        if (axi_master==CHIP) mig_rvalid_cnt <= mig_rvalid_cnt + 32'd1;
                    end
                end
            endcase
        end
    end


    //************************************************************
    // Self wstrb generation 
    //************************************************************

    always @(*) begin
        if (wcnt == 8'd0) begin
            if (wstart && s_axi_wready && s_axi_wvalid && chip_store_byte4) s_axi_wstrb = 32'h0000_000f << s_axi_awaddr[4:0];
            else if (chip_store_byte4_buf) s_axi_wstrb = 32'h0000_000f << awaddr_buf[4:0];
            else                           s_axi_wstrb = 32'hffff_ffff << awaddr_buf[4:0];
        end
        else s_axi_wstrb = 32'hffff_ffff;
    end

    always @(posedge clk or negedge rstn) begin
        if (~rstn) begin
            chip_store_byte4_buf <= 1'b0;
        end
        else begin
            // capture chip_store_byte4
            if (wstart) begin
                chip_store_byte4_buf <= chip_store_byte4;
            end
            else begin
                chip_store_byte4_buf <= 1'b0;
            end
        end
    end



    //************************************************************
    // Instantiate MIG module
    //************************************************************

    always @(posedge clk) begin
        aresetn <= ~rst;
    end

    xem7360_k160t_mig u_xem7360_k160t_mig
    (
        // Memory interface ports
        .ddr3_addr                      (ddr3_addr              ),
        .ddr3_ba                        (ddr3_ba                ),
        .ddr3_cas_n                     (ddr3_cas_n             ),
        .ddr3_ck_n                      (ddr3_ck_n              ),
        .ddr3_ck_p                      (ddr3_ck_p              ),
        .ddr3_cke                       (ddr3_cke               ),
        .ddr3_ras_n                     (ddr3_ras_n             ),
        .ddr3_we_n                      (ddr3_we_n              ),
        .ddr3_dq                        (ddr3_dq                ),
        .ddr3_dqs_n                     (ddr3_dqs_n             ),
        .ddr3_dqs_p                     (ddr3_dqs_p             ),
        .ddr3_reset_n                   (ddr3_reset_n           ),
        .init_calib_complete            (init_calib_complete    ),
        .ddr3_cs_n                      (ddr3_cs_n              ),
        .ddr3_dm                        (ddr3_dm                ),
        .ddr3_odt                       (ddr3_odt               ),

        // Application interface ports
        .ui_clk                         (clk                    ),  // output
        .ui_clk_sync_rst                (rst                    ),  // output
        .mmcm_locked                    (mmcm_locked            ),  // not used
        .aresetn                        (aresetn                ),
        .app_sr_req                     (1'b0                   ),
        .app_ref_req                    (1'b0                   ),
        .app_zq_req                     (1'b0                   ),
        .app_sr_active                  (                       ),
        .app_ref_ack                    (                       ),
        .app_zq_ack                     (                       ),

        // Slave Interface Write Address Ports
        .s_axi_awid                     (1'b0                   ),
        .s_axi_awaddr                   ({3'b0, s_axi_awaddr}   ),
        .s_axi_awlen                    (s_axi_awlen            ),
        .s_axi_awsize                   (3'b101                 ),
        .s_axi_awburst                  (2'b01                  ),
        .s_axi_awlock                   (1'b0                   ),
        .s_axi_awcache                  (4'b0                   ),
        .s_axi_awprot                   (3'b010                 ),
        .s_axi_awqos                    (4'h0                   ),
        .s_axi_awvalid                  (s_axi_awvalid          ),
        .s_axi_awready                  (s_axi_awready          ),

        // Slave Interface Write Data Ports
        .s_axi_wdata                    (s_axi_wdata            ),
        .s_axi_wstrb                    (s_axi_wstrb            ),
        .s_axi_wlast                    (s_axi_wlast            ),
        .s_axi_wvalid                   (s_axi_wvalid           ),
        .s_axi_wready                   (s_axi_wready           ),

        // Slave Interface Write Response Ports
        .s_axi_bid                      (s_axi_bid              ),
        .s_axi_bresp                    (s_axi_bresp            ),
        .s_axi_bvalid                   (s_axi_bvalid           ),
        .s_axi_bready                   (1'b1                   ),

        // Slave Interface Read Address Ports
        .s_axi_arid                     (1'b0                   ),
        .s_axi_araddr                   ({3'b0, s_axi_araddr}   ),
        .s_axi_arlen                    (s_axi_arlen            ),
        .s_axi_arsize                   (3'b101                 ),
        .s_axi_arburst                  (2'b01                  ),
        .s_axi_arlock                   (1'b0                   ),
        .s_axi_arcache                  (4'b0                   ),
        .s_axi_arprot                   (3'b010                 ),
        .s_axi_arqos                    (4'h0                   ),
        .s_axi_arvalid                  (s_axi_arvalid          ),
        .s_axi_arready                  (s_axi_arready          ),

        // Slave Interface Read Data Ports
        .s_axi_rid                      (s_axi_rid              ),
        .s_axi_rdata                    (s_axi_rdata            ),
        .s_axi_rresp                    (s_axi_rresp            ),
        .s_axi_rlast                    (s_axi_rlast            ),
        .s_axi_rvalid                   (s_axi_rvalid           ),
        .s_axi_rready                   (s_axi_rready           ),

        // System Clock Ports
        .sys_clk_p                      (sys_clk_p              ),
        .sys_clk_n                      (sys_clk_n              ),
        .device_temp                    (                       ),

        .sys_rst                        (~okRstn                )    // active-high
    );



endmodule