//`define SKIP_CALIB 1
// `define LOOPBACK_TEST 1
// `define CLK_EXT 1   // use external clock, comment out this line to generate clk internally and use this for chip
`define BUILTIN_FIFO 1
// `define DEBUG_FIFO 1