//////////////////////////////////////////////////////////////////////////////////
// Engineer: Kim Beomseok
// Contact: kimbss470@snu.ac.kr
// 
// Create Date: 15/07/2024 
// Design Name: OpalKelly frontpanel for USB3 in Verilog
// Module Name: okFrontPanel
// Project Name: 2024TapeOut
// Target Devices: XEM7360-K160T
// Tool versions: 2024.1
// Description: 
//
//////////////////////////////////////////////////////////////////////////////////

module okFrontPanel (
    input  wire          init_calib_done,
    input  wire          rstn, // generated by clock wizard 

    output wire          okClk,
    input  wire [  4:0]  okUH,
    output wire [  2:0]  okHU,
    inout  wire [ 31:0]  okUHU,
    inout  wire          okAA,
    output wire          okRstn,   // input to clock wizard and MIG


    /* okFP <-> Chip */
    input  wire          chip_clk,
    output wire          chip_network_start,
    output wire          chip_single_rate,
    output wire [  5:0]  chip_n_layers,
    output wire          chip_infinite_loop,
    output wire [ 15:0]  wait_chip_cnt,
    input  wire          chip_network_done,
    input  wire [31:0]   chip_done_network_cnt,
    input  wire          chip_layer_done,    // buffered for done from chip, synchronized with clk_for_chip_out
    input  wire [ 30:0]  chip_clk_cnt,


    /* AXI-interface (okFP <-> MIG ) */
    input  wire          mig_clk,
    output reg           mig_abort,
    output reg           axi_master,
    output wire [ 27:0]  axi_awaddr,     // Write address
    output wire [  7:0]  axi_awlen,
    output wire          axi_awvalid,
    input  wire          axi_awready,

    output wire [255:0]  axi_wdata,      // Write data 
    output wire          axi_wvalid,
    input  wire          axi_wready,

    output wire [ 27:0]  axi_araddr,     // Read address
    output wire [  7:0]  axi_arlen,
    output wire          axi_arvalid,
    input  wire          axi_arready,

    input  wire [255:0]  axi_rdata,      // Read data
    input  wire          axi_rvalid,
    output wire          axi_rready,

    /* Debug (ChipInterface) */
    input  wire [  7:0]  start_cnt,
    input  wire [  7:0]  done_cnt,
    input  wire [ 31:0]  arvalid_cnt,
    input  wire [  7:0]  arready_cnt,
    input  wire [ 31:0]  rvalid_cnt,
    input  wire [ 31:0]  awvalid_cnt,
    input  wire [  7:0]  awready_cnt,
    input  wire [ 31:0]  wvalid_cnt,
    input  wire [ 27:0]  araddr_hist [0:63],
    input  wire [  7:0]  arlen_hist  [0:63],
    input  wire [255:0]  rdata_hist  [0:63],
    input  wire [ 27:0]  awaddr_hist [0:63],
    input  wire [  7:0]  awlen_hist  [0:63],
    // output wire [255:0]  wdata_hist  [0:255]

    input  wire [  3:0]  ttf_axvalid,

    /* FIFO for cycle level debugging of fpga2chip signals */
    output wire          debug_fifo_fpga2chip_read,
    input  wire          debug_fifo_fpga2chip_rd_en,
    output wire          pipe_out_ready_debug_fpga2chip,
    input  wire          pipe_out_valid_debug_fpga2chip,
    input  wire [ 31:0]  pipe_dout_debug_fpga2chip,

    /* FIFO for cycle level debugging of chip2fpga signals */
    output wire          debug_fifo_chip2fpga_read,
    input  wire          debug_fifo_chip2fpga_rd_en,
    output wire          pipe_out_ready_debug_chip2fpga,
    input  wire          pipe_out_valid_debug_chip2fpga,
    input  wire [ 31:0]  pipe_dout_debug_chip2fpga,

    /* FIFO for axaddr and axlen handshaking debugging */
    output wire          debug_fifo_axaddr_read,
    input  wire          debug_fifo_axaddr_rd_en,
    output wire          pipe_out_ready_debug_axaddr,
    input  wire          pipe_out_valid_debug_axaddr,
    input  wire [ 31:0]  pipe_dout_debug_axaddr,

    /* FIFO for rdata transfer debugging */
    output wire          debug_fifo_rdata_read,
    input  wire          debug_fifo_rdata_rd_en,
    output wire          pipe_out_ready_debug_rdata,
    input  wire          pipe_out_valid_debug_rdata,
    input  wire [ 31:0]  pipe_dout_debug_rdata,

    /* FIFO for wdata transfer debugging */
    output wire          debug_fifo_wdata_read,
    input  wire          debug_fifo_wdata_rd_en,
    output wire          pipe_out_ready_debug_wdata,
    input  wire          pipe_out_valid_debug_wdata,
    input  wire [ 31:0]  pipe_dout_debug_wdata,


    /* Debug of regular FIFOs btw chip <-> MIG */
    input  wire          araddr_fifo_rd_en_debug,
    input  wire          araddr_fifo_wr_en_debug,
    input  wire          araddr_fifo_valid_debug, 
    input  wire          araddr_fifo_empty_debug, 
    input  wire          araddr_fifo_full_debug, 
    input  wire          araddr_fifo_prog_full_debug, 
 
    input  wire          awaddr_fifo_rd_en_debug,
    input  wire          awaddr_fifo_wr_en_debug,
    input  wire          awaddr_fifo_valid_debug, 
    input  wire          awaddr_fifo_empty_debug, 
    input  wire          awaddr_fifo_full_debug, 
    input  wire          awaddr_fifo_prog_full_debug, 
 
    input  wire          rdata_fifo_rd_en_debug,
    input  wire          rdata_fifo_wr_en_debug,
    input  wire          rdata_fifo_valid_debug, 
    input  wire          rdata_fifo_empty_debug, 
    input  wire          rdata_fifo_full_debug, 
    input  wire          rdata_fifo_prog_full_debug, 
 
    input  wire          wdata_fifo_rd_en_debug,
    input  wire          wdata_fifo_wr_en_debug,
    input  wire          wdata_fifo_valid_debug, 
    input  wire          wdata_fifo_empty_debug, 
    input  wire          wdata_fifo_full_debug, 
    input  wire          wdata_fifo_prog_full_debug,

    /* Debug (DDR3Interface) */
    input  wire          s_axi_arready_debug,
    input  wire          s_axi_rvalid_debug,
    input  wire          s_axi_wstate_debug,
    input  wire          s_axi_wready_debug,
    input  wire [ 31:0]  mig_rstate_cnt,
    input  wire [ 31:0]  mig_rvalid_cnt,
    input  wire [ 31:0]  mig_wstate_cnt,
    input  wire [ 31:0]  mig_wvalid_cnt
);
    `include "params.vh"
    localparam NUM_EP_OUT = 30;

    // states
    localparam S_IDLE                = 4'd0;
    localparam S_DRAM_WRITE          = 4'd1;
    localparam S_DRAM_READ           = 4'd2;
    localparam S_EXECUTE_NET         = 4'd3;
    localparam S_FIFO_FPGA2CHIP_READ = 4'd4;
    localparam S_FIFO_CHIP2FPGA_READ = 4'd5;
    localparam S_FIFO_AXADDR_READ    = 4'd6;
    localparam S_FIFO_RDATA_READ     = 4'd7;
    localparam S_FIFO_WDATA_READ     = 4'd8;

    // cmd 
    localparam CMD_DRAM_WRITE          = 32'b000000001;
    localparam CMD_DRAM_READ           = 32'b000000010;
    localparam CMD_EXECUTE_NET         = 32'b000000100;
    localparam CMD_FIFO_FPGA2CHIP_READ = 32'b000001000;
    localparam CMD_FIFO_CHIP2FPGA_READ = 32'b000010000;
    localparam CMD_FIFO_AXADDR_READ    = 32'b000100000;
    localparam CMD_FIFO_RDATA_READ     = 32'b001000000;
    localparam CMD_FIFO_WDATA_READ     = 32'b010000000;
    localparam CMD_ABORT               = 32'b100000000;

    // AXI-master
    localparam OKFP = 1'd0;
    localparam CHIP = 1'd1;

    // FIFO
    localparam FIFO_HEADROOM = 20;

    //************************************************************
    //  Wires & Regs 
    //************************************************************

    /* Target interface bus */
    // wire                     okClk;
    wire [112:0]             okHE;
    wire [64:0]              okEH;
    wire [65*NUM_EP_OUT-1:0] okEHx;

    /* Endpoint connections */
    wire [31:0]  ep00wire;    // <-- rstn
    wire [31:0]  ep01wire;    // <-- addr
    wire [31:0]  ep02wire;    // <-- len (bytes)
    wire [31:0]  ep03wire;    // <-- single/dual-rate (chip supports only single-rate..)
    wire [31:0]  ep04wire;    // <-- n_layers
    wire [31:0]  ep07wire;    // <-- infinite loop mode
    wire [31:0]  ep08wire;    // <-- wait_chip_cnt
    wire [31:0]  ep20wire;    // --> current_state
    wire [31:0]  ep21wire;    // --> clk_cnt

    wire [31:0]  ep05wire;    // for debug
    wire [31:0]  ep06wire;    // for debug
    wire [31:0]  ep22wire;    // for debug
    wire [31:0]  ep23wire;    // for debug
    wire [31:0]  ep24wire;    // for debug
    wire [31:0]  ep25wire;    // for debug
    wire [31:0]  ep26wire;    // for debug
    wire [31:0]  ep27wire;    // for debug
    wire [31:0]  ep28wire;    // for debug
    wire [31:0]  ep29wire;    // for debug
    wire [31:0]  ep30wire;    // for debug
    wire [31:0]  ep31wire;    // for debug
    wire [31:0]  ep32wire;    // for debug
    wire [31:0]  ep33wire;    // for debug
    wire [31:0]  ep34wire;    // for debug
    wire [31:0]  ep35wire;    // for debug
    wire [31:0]  ep36wire;    // for debug
    wire [31:0]  ep37wire;    // for debug
    wire [31:0]  ep38wire;    // for debug
    wire [31:0]  ep39wire;    // for debug

    wire [31:0]  ep40trig;    // <-- cmd
    wire [31:0]  ep60trig;    // --> init_calib_done
    wire [31:0]  ep61trig;    // --> network_done
    wire [31:0]  ep62trig;    // --> layer_done

    wire         pipe_in_ready;
    wire         pipe_in_valid;
    wire [31:0]  pipe_din;
    wire         pipe_out_ready;
    reg          pipe_out_ready_buf;
    wire         pipe_out_valid;
    wire [31:0]  pipe_dout;


    /*  Reordering axi data  */ 
    wire [255:0] axi_wdata_pre_ord;
    wire [255:0] axi_rdata_aft_ord;


    /*  FIFOs between okFP <-> MIG  */ 
    wire         fifo_rst;
    wire         araddr_fifo_wr_en; 
    wire         araddr_fifo_rd_en; 
    wire [35:0]  araddr_fifo_din; 
    wire [35:0]  araddr_fifo_dout; 
    wire         araddr_fifo_valid; 
    wire         araddr_fifo_empty; 
    wire         araddr_fifo_full; 
    wire         araddr_fifo_prog_full; 

    wire         awaddr_fifo_wr_en; 
    wire         awaddr_fifo_rd_en; 
    wire [35:0]  awaddr_fifo_din; 
    wire [35:0]  awaddr_fifo_dout; 
    wire         awaddr_fifo_valid; 
    wire         awaddr_fifo_empty; 
    wire         awaddr_fifo_full; 
    wire         awaddr_fifo_prog_full; 

    wire         rdata_fifo_wr_en; 
    wire         rdata_fifo_rd_en; 
    wire [255:0] rdata_fifo_din; 
    wire [ 31:0] rdata_fifo_dout; 
    wire         rdata_fifo_valid; 
    wire         rdata_fifo_empty; 
    wire         rdata_fifo_full; 
    wire         rdata_fifo_prog_full; 

    wire         wdata_fifo_wr_en; 
    wire         wdata_fifo_rd_en; 
    wire [ 31:0] wdata_fifo_din; 
    wire [255:0] wdata_fifo_dout; 
    wire         wdata_fifo_valid; 
    wire         wdata_fifo_empty; 
    wire         wdata_fifo_full; 
    wire         wdata_fifo_prog_full; 


    /*  FIFOs between okFP <-> chip */ 
    wire         ok2chip_fifo_wr_en;
    wire         ok2chip_fifo_rd_en;
    wire [7:0]   ok2chip_fifo_din;
    wire [7:0]   ok2chip_fifo_dout;
    wire         ok2chip_fifo_valid;
    wire         ok2chip_fifo_empty;
    wire         ok2chip_fifo_full;
    wire         ok2chip_fifo_prog_full;

    wire         chip2ok_fifo_wr_en;
    wire         chip2ok_fifo_rd_en;
    wire [31:0]  chip2ok_fifo_din;
    wire [31:0]  chip2ok_fifo_dout;
    wire         chip2ok_fifo_valid;
    wire         chip2ok_fifo_empty;
    wire         chip2ok_fifo_full;
    wire         chip2ok_fifo_prog_full;

    /* okFP -> Chip signals  */ 
    
    
    /* FSM */
    reg  [3:0]   state;

    wire [31:0]  cmd;
    reg  [31:0]  cmd_buf;
    wire         abort;
    wire         dram_write_done;
    wire         dram_read_done;
    reg  [11:0]  i_transfer;
    reg  [13:0]  len;    // bytes
    reg  [27:0]  addr;
    wire [7:0]   axi_axlen;
    reg          network_start;
    reg          single_rate;
    reg  [5:0]   n_layers;
    reg          infinite_loop;
    
    wire         network_done;
    reg          network_done_buf;
    reg          layer_done_buf0;   // synchronizer
    reg          layer_done_buf1;   // synchronizer
    wire [30:0]  clk_cnt;
    reg  [30:0]  clk_cnt_buf;

    wire         debug_fifo_fpga2chip_read_done;
    wire         debug_fifo_chip2fpga_read_done;
    wire         debug_fifo_axaddr_read_done;
    wire         debug_fifo_rdata_read_done;
    wire         debug_fifo_wdata_read_done;
    


    //************************************************************
    // Instantiate the okHost and connect endpoints
    //************************************************************

    /* okHost */
    okHost okHI(
        .okUH (okUH),
        .okHU (okHU),
        .okUHU(okUHU),
        .okAA (okAA),
        .okClk(okClk),
        .okHE (okHE),
        .okEH (okEH)
    );

    /* okWireOR */
    okWireOR #(.N(NUM_EP_OUT)) wireOR (.okEH(okEH), .okEHx(okEHx));

    /* okWireIn */
    okWireIn  wireIn00 (.okHE(okHE), .ep_addr(8'h00), .ep_dataout(ep00wire));    // rstn
    okWireIn  wireIn01 (.okHE(okHE), .ep_addr(8'h01), .ep_dataout(ep01wire));    // addr
    okWireIn  wireIn02 (.okHE(okHE), .ep_addr(8'h02), .ep_dataout(ep02wire));    // len
    okWireIn  wireIn03 (.okHE(okHE), .ep_addr(8'h03), .ep_dataout(ep03wire));    // single-rate 
    okWireIn  wireIn04 (.okHE(okHE), .ep_addr(8'h04), .ep_dataout(ep04wire));    // n_layers 
    okWireIn  wireIn05 (.okHE(okHE), .ep_addr(8'h05), .ep_dataout(ep05wire));    // (DEBUG) read_or_write, 0 for read 1 for write
    okWireIn  wireIn06 (.okHE(okHE), .ep_addr(8'h06), .ep_dataout(ep06wire));    // (DEBUG) history idx
    okWireIn  wireIn07 (.okHE(okHE), .ep_addr(8'h07), .ep_dataout(ep07wire));    // infinite loop mode
    okWireIn  wireIn08 (.okHE(okHE), .ep_addr(8'h08), .ep_dataout(ep08wire));    // wait_chip_cnt


    /* okWireOut */
    okWireOut wireOut20 (.okHE(okHE), .okEH(okEHx[ 0*65 +: 65]), .ep_addr(8'h20), .ep_datain(ep20wire));    // current state
    okWireOut wireOut21 (.okHE(okHE), .okEH(okEHx[ 1*65 +: 65]), .ep_addr(8'h21), .ep_datain(ep21wire));    // clk_cnt_buf
    okWireOut wireOut22 (.okHE(okHE), .okEH(okEHx[ 2*65 +: 65]), .ep_addr(8'h22), .ep_datain(ep22wire));    // (DEBUG) chip_clk_cnt
    okWireOut wireOut23 (.okHE(okHE), .okEH(okEHx[ 3*65 +: 65]), .ep_addr(8'h23), .ep_datain(ep23wire));    // (DEBUG) chip_done_network_cnt
    okWireOut wireOut24 (.okHE(okHE), .okEH(okEHx[ 4*65 +: 65]), .ep_addr(8'h24), .ep_datain(ep24wire));    // (DEBUG) axaddr_hist[hist_idx]
    okWireOut wireOut25 (.okHE(okHE), .okEH(okEHx[ 5*65 +: 65]), .ep_addr(8'h25), .ep_datain(ep25wire));    // (DEUBG) axlen_hist[hist_idx]
    okWireOut wireOut26 (.okHE(okHE), .okEH(okEHx[ 6*65 +: 65]), .ep_addr(8'h26), .ep_datain(ep26wire));    // (DEBUG) rdata_hist[hist_idx][32*7+:32] -> arvalid_cnt
    okWireOut wireOut27 (.okHE(okHE), .okEH(okEHx[ 7*65 +: 65]), .ep_addr(8'h27), .ep_datain(ep27wire));    // (DEBUG) rdata_hist[hist_idx][32*6+:32] -> rvalid_cnt
    okWireOut wireOut28 (.okHE(okHE), .okEH(okEHx[ 8*65 +: 65]), .ep_addr(8'h28), .ep_datain(ep28wire));    // (DEBUG) rdata_hist[hist_idx][32*5+:32] -> awvalid_cnt
    okWireOut wireOut29 (.okHE(okHE), .okEH(okEHx[ 9*65 +: 65]), .ep_addr(8'h29), .ep_datain(ep29wire));    // (DEBUG) rdata_hist[hist_idx][32*4+:32] -> wvalid_cnt
    okWireOut wireOut30 (.okHE(okHE), .okEH(okEHx[10*65 +: 65]), .ep_addr(8'h30), .ep_datain(ep30wire));    // (DEBUG) rdata_hist[hist_idx][32*3+:32] -> mig_rstate_cnt
    okWireOut wireOut31 (.okHE(okHE), .okEH(okEHx[11*65 +: 65]), .ep_addr(8'h31), .ep_datain(ep31wire));    // (DEBUG) rdata_hist[hist_idx][32*2+:32] -> mig_rvalid_cnt
    okWireOut wireOut32 (.okHE(okHE), .okEH(okEHx[12*65 +: 65]), .ep_addr(8'h32), .ep_datain(ep32wire));    // (DEBUG) rdata_hist[hist_idx][32*1+:32] -> mig_wstate_cnt
    okWireOut wireOut33 (.okHE(okHE), .okEH(okEHx[13*65 +: 65]), .ep_addr(8'h33), .ep_datain(ep33wire));    // (DEBUG) rdata_hist[hist_idx][32*0+:32] -> mig_wvalid_cnt
    okWireOut wireOut34 (.okHE(okHE), .okEH(okEHx[14*65 +: 65]), .ep_addr(8'h34), .ep_datain(ep34wire));    // (DEBUG) DDR3Interface wstate, wready, rstate, rready
    okWireOut wireOut35 (.okHE(okHE), .okEH(okEHx[15*65 +: 65]), .ep_addr(8'h35), .ep_datain(ep35wire));    // (DEBUG) {mig wstate_cnt, rstate_cnt}
    okWireOut wireOut36 (.okHE(okHE), .okEH(okEHx[16*65 +: 65]), .ep_addr(8'h36), .ep_datain(ep36wire));    // (DEBUG) chip<=>mig fifo status
    okWireOut wireOut37 (.okHE(okHE), .okEH(okEHx[17*65 +: 65]), .ep_addr(8'h37), .ep_datain(ep37wire));    // (DEBUG) ttf_axvalid
    okWireOut wireOut38 (.okHE(okHE), .okEH(okEHx[18*65 +: 65]), .ep_addr(8'h38), .ep_datain(ep38wire));    // (DEBUG) {awvalid_cnt, wvalid_cnt}
    okWireOut wireOut39 (.okHE(okHE), .okEH(okEHx[19*65 +: 65]), .ep_addr(8'h39), .ep_datain(ep39wire));    // (DEBUG) {debug_chip_network_done_cnt, debug_ok_network_done_cnt}

    /* okTriggerIn */
    okTriggerIn  trigIn40 (.okHE(okHE), .ep_addr(8'h40), .ep_clk(okClk), .ep_trigger(ep40trig));     // cmd (start)

    /* okTriggerOut */
    okTriggerOut trigOut60 (.okHE(okHE), .okEH(okEHx[20*65 +: 65]), .ep_addr(8'h60), .ep_clk(okClk), .ep_trigger(ep60trig));    // init_calib_done 
    okTriggerOut trigOut61 (.okHE(okHE), .okEH(okEHx[21*65 +: 65]), .ep_addr(8'h61), .ep_clk(okClk), .ep_trigger(ep61trig));    // network_done
    okTriggerOut trigOut62 (.okHE(okHE), .okEH(okEHx[22*65 +: 65]), .ep_addr(8'h62), .ep_clk(okClk), .ep_trigger(ep62trig));    // layer_done (optional)
    
    /* okBTPipeIn */
    okBTPipeIn  btPipeIn  (.okHE(okHE), .okEH(okEHx[23*65 +:65]), .ep_addr(8'h80), .ep_dataout(pipe_din), .ep_write(pipe_in_valid), .ep_blockstrobe(), .ep_ready(pipe_in_ready));

    /* okBTPipeOut */
    okBTPipeOut btPipeOutA0 (.okHE(okHE), .okEH(okEHx[24*65 +:65]), .ep_addr(8'hA0), .ep_datain(pipe_dout), .ep_read(pipe_out_ready), .ep_blockstrobe(), .ep_ready(pipe_out_valid));
    okBTPipeOut btPipeOutA1 (.okHE(okHE), .okEH(okEHx[25*65 +:65]), .ep_addr(8'hA1), .ep_datain(pipe_dout_debug_fpga2chip), .ep_read(pipe_out_ready_debug_fpga2chip), .ep_blockstrobe(), .ep_ready(pipe_out_valid_debug_fpga2chip));
    okBTPipeOut btPipeOutA2 (.okHE(okHE), .okEH(okEHx[26*65 +:65]), .ep_addr(8'hA2), .ep_datain(pipe_dout_debug_chip2fpga), .ep_read(pipe_out_ready_debug_chip2fpga), .ep_blockstrobe(), .ep_ready(pipe_out_valid_debug_chip2fpga));
    okBTPipeOut btPipeOutA3 (.okHE(okHE), .okEH(okEHx[27*65 +:65]), .ep_addr(8'hA3), .ep_datain(pipe_dout_debug_axaddr), .ep_read(pipe_out_ready_debug_axaddr), .ep_blockstrobe(), .ep_ready(pipe_out_valid_debug_axaddr));
    okBTPipeOut btPipeOutA4 (.okHE(okHE), .okEH(okEHx[28*65 +:65]), .ep_addr(8'hA4), .ep_datain(pipe_dout_debug_rdata), .ep_read(pipe_out_ready_debug_rdata), .ep_blockstrobe(), .ep_ready(pipe_out_valid_debug_rdata));
    okBTPipeOut btPipeOutA5 (.okHE(okHE), .okEH(okEHx[29*65 +:65]), .ep_addr(8'hA5), .ep_datain(pipe_dout_debug_wdata), .ep_read(pipe_out_ready_debug_wdata), .ep_blockstrobe(), .ep_ready(pipe_out_valid_debug_wdata));



    //************************************************************
    // Endpoint Wire Connections
    //************************************************************

    assign okRstn   = ~ep00wire[0];    // active-low

    assign wait_chip_cnt = ep08wire[15:0];
    assign ep20wire = {28'd0, state};
    assign ep21wire = {1'b0, clk_cnt_buf};
    assign ep22wire = {1'b0, chip_clk_cnt};   // (chip-clk domain) not buffered -> used only for infinite loop mode
    assign ep23wire = chip_done_network_cnt;  // (chip-clk domain) used only for infinite loop mode

    assign cmd      = ep40trig;
    assign ep60trig = {31'd0, init_calib_done};
    assign ep61trig = {31'b0, network_done_buf};
    assign ep62trig = {31'b0, layer_done_buf1};   

    always @(posedge okClk) begin
        layer_done_buf0 <= chip_layer_done;
        layer_done_buf1 <= layer_done_buf0; 
    end


    //************************************************************
    // DRAM Read/Write FSM
    //************************************************************

    assign axi_axlen                       = len[13:5] - 9'd1;    // 32bytes per each transfer
    assign dram_write_done                 = (state == S_DRAM_WRITE) && (len[13:2] == i_transfer);
    assign dram_read_done                  = (state == S_DRAM_READ ) && (len[13:2] == i_transfer);
    assign debug_fifo_fpga2chip_read       = (state == S_FIFO_FPGA2CHIP_READ);
    assign debug_fifo_chip2fpga_read       = (state == S_FIFO_CHIP2FPGA_READ);
    assign debug_fifo_axaddr_read          = (state == S_FIFO_AXADDR_READ   );
    assign debug_fifo_rdata_read           = (state == S_FIFO_RDATA_READ    );
    assign debug_fifo_wdata_read           = (state == S_FIFO_WDATA_READ    );
    assign debug_fifo_fpga2chip_read_done  = (state == S_FIFO_FPGA2CHIP_READ) && (len[13:2] == i_transfer);
    assign debug_fifo_chip2fpga_read_done  = (state == S_FIFO_CHIP2FPGA_READ) && (len[13:2] == i_transfer);
    assign debug_fifo_axaddr_read_done     = (state == S_FIFO_AXADDR_READ   ) && (len[13:2] == i_transfer);
    assign debug_fifo_rdata_read_done      = (state == S_FIFO_RDATA_READ    ) && (len[13:2] == i_transfer);
    assign debug_fifo_wdata_read_done      = (state == S_FIFO_WDATA_READ    ) && (len[13:2] == i_transfer);

    assign abort = (cmd == CMD_ABORT);

    always @(posedge okClk or negedge rstn) begin
        if (~rstn) begin
            state  <= S_IDLE;
        end
        else begin
            case (state)
                S_IDLE: begin
                    if      (cmd == CMD_DRAM_WRITE         ) state <= S_DRAM_WRITE;
                    else if (cmd == CMD_DRAM_READ          ) state <= S_DRAM_READ;
                    else if (cmd == CMD_EXECUTE_NET        ) state <= S_EXECUTE_NET;
                    else if (cmd == CMD_FIFO_FPGA2CHIP_READ) state <= S_FIFO_FPGA2CHIP_READ;
                    else if (cmd == CMD_FIFO_CHIP2FPGA_READ) state <= S_FIFO_CHIP2FPGA_READ;
                    else if (cmd == CMD_FIFO_AXADDR_READ   ) state <= S_FIFO_AXADDR_READ;
                    else if (cmd == CMD_FIFO_RDATA_READ    ) state <= S_FIFO_RDATA_READ;
                    else if (cmd == CMD_FIFO_WDATA_READ    ) state <= S_FIFO_WDATA_READ;
                    else                                     state <= S_IDLE;
                end
                S_DRAM_WRITE: begin
                    if (dram_write_done) state <= S_IDLE;
                end
                S_DRAM_READ: begin
                    if (dram_read_done) state <= S_IDLE;
                end
                S_EXECUTE_NET: begin
                    if (abort || network_done) state <= S_IDLE;
                end
                S_FIFO_FPGA2CHIP_READ: begin
                    if (abort || debug_fifo_fpga2chip_read_done) state <= S_IDLE;
                end
                S_FIFO_CHIP2FPGA_READ: begin
                    if (abort || debug_fifo_chip2fpga_read_done) state <= S_IDLE;
                end
                S_FIFO_AXADDR_READ: begin
                    if (abort || debug_fifo_axaddr_read_done) state <= S_IDLE;
                end
                S_FIFO_RDATA_READ: begin
                    if (abort || debug_fifo_rdata_read_done) state <= S_IDLE;
                end
                S_FIFO_WDATA_READ: begin
                    if (abort || debug_fifo_wdata_read_done) state <= S_IDLE;
                end
            endcase
        end
    end

    always @(posedge okClk or negedge rstn) begin
        if (~rstn) begin
            cmd_buf          <= 'd0;
            addr             <= 'd0;
            len              <= 'd0;
            axi_master       <= OKFP;
            i_transfer       <= 12'd0;

            network_start    <= 1'b0;
            network_done_buf <= 1'b0;
            single_rate      <= 1'b0;
            n_layers         <= 6'd0;
            infinite_loop    <= 1'b0;
            clk_cnt_buf      <= 31'd0;
        end
        else begin
            
            cmd_buf <= cmd;

            case (state)
                S_IDLE: begin
                    if ((cmd == CMD_DRAM_WRITE) || (cmd == CMD_DRAM_READ)) begin
                        addr <= ep01wire[27:0];   // dram addr
                        len  <= ep02wire[13:0];   // bytes to write/read
                    end
                    else if ((cmd == CMD_FIFO_FPGA2CHIP_READ) || (cmd == CMD_FIFO_CHIP2FPGA_READ) 
                            || (cmd == CMD_FIFO_AXADDR_READ) || (cmd == CMD_FIFO_RDATA_READ) 
                            || (cmd == CMD_FIFO_WDATA_READ)) begin
                        addr <= 'd0;
                        len  <= ep02wire[13:0];    // byte to read  
                    end
                    else begin
                        addr <= 'd0;
                        len  <= 'd0;
                    end

                    if (cmd == CMD_EXECUTE_NET) axi_master <= CHIP;
                    else                        axi_master <= OKFP;

                    i_transfer       <= 12'd0;

                    if (cmd == CMD_EXECUTE_NET) begin
                        network_start <= 1'b1;
                        single_rate   <= ep03wire[0];
                        n_layers      <= ep04wire[5:0];
                        infinite_loop <= ep07wire[0];
                    end
                    else begin
                        network_start <= 1'b0;
                        single_rate   <= 1'b0;
                        n_layers      <= 6'd0;
                        infinite_loop <= 1'b0;
                    end

                    network_done_buf <= 1'b0;
                    // clk_cnt_buf      <= 31'd0;
                end

                S_DRAM_WRITE: begin
                    if (dram_write_done) begin
                        i_transfer <= 12'd0;
                    end
                    else if (pipe_in_valid) begin
                        i_transfer <= i_transfer + 12'd1;
                    end
                end

                S_DRAM_READ: begin
                    if (dram_read_done) begin
                        i_transfer <= 12'd0;
                    end
                    else if (rdata_fifo_rd_en) begin
                        i_transfer <= i_transfer + 12'd1;
                    end
                end

                S_EXECUTE_NET: begin
                    network_start <= 1'b0;
                    network_done_buf <= network_done;
                    if (network_done) begin
                        // Set triggerOut
                        clk_cnt_buf      <= clk_cnt;
                    end
                end

                S_FIFO_FPGA2CHIP_READ: begin
                    if (debug_fifo_fpga2chip_read_done) begin
                        i_transfer <= 12'd0;
                    end
                    else if (debug_fifo_fpga2chip_rd_en) begin
                        i_transfer <= i_transfer + 12'd1;
                    end
                end

                S_FIFO_CHIP2FPGA_READ: begin
                    if (debug_fifo_chip2fpga_read_done) begin
                        i_transfer <= 12'd0;
                    end
                    else if (debug_fifo_chip2fpga_rd_en) begin
                        i_transfer <= i_transfer + 12'd1;
                    end
                end

                S_FIFO_AXADDR_READ: begin
                    if (debug_fifo_axaddr_read_done) begin
                        i_transfer <= 12'd0;
                    end
                    else if (debug_fifo_axaddr_rd_en) begin
                        i_transfer <= i_transfer + 12'd1;
                    end
                end

                S_FIFO_RDATA_READ: begin
                    if (debug_fifo_rdata_read_done) begin
                        i_transfer <= 12'd0;
                    end
                    else if (debug_fifo_rdata_rd_en) begin
                        i_transfer <= i_transfer + 12'd1;
                    end
                end
                
                S_FIFO_WDATA_READ: begin
                    if (debug_fifo_wdata_read_done) begin
                        i_transfer <= 12'd0;
                    end
                    else if (debug_fifo_wdata_rd_en) begin
                        i_transfer <= i_transfer + 12'd1;
                    end
                end
            endcase
        end
    end



    //************************************************************
    // Instantiate FIFOs between okFP <-> MIG
    //************************************************************

    assign fifo_rst = ~rstn;    // active-high

    /* awaddr fifo (okFP -> MIG) */
    awaddr_fifo_36_128 awaddr_fifo (
        .rst                (fifo_rst              ),    // active-high
        .wr_clk             (okClk                 ),
        .rd_clk             (mig_clk               ),
        .din                (awaddr_fifo_din       ),
        .wr_en              (awaddr_fifo_wr_en     ),
        .rd_en              (awaddr_fifo_rd_en     ),
        .dout               (awaddr_fifo_dout      ),
        .full               (awaddr_fifo_full      ),
        .empty              (awaddr_fifo_empty     ),
        .valid              (awaddr_fifo_valid     ),
        .prog_full_thresh   (7'd127-FIFO_HEADROOM  ),
        .prog_full          (awaddr_fifo_prog_full )
    );

    /* wdata fifo (okFP -> MIG) */
    wdata_fifo_w32_1024_r256_128 wdata_fifo (
        .rst                (fifo_rst              ),    // active-high
        .wr_clk             (okClk                 ),
        .rd_clk             (mig_clk               ),
        .din                (wdata_fifo_din        ),
        .wr_en              (wdata_fifo_wr_en      ),
        .rd_en              (wdata_fifo_rd_en      ),
        .dout               (wdata_fifo_dout       ),
        .full               (wdata_fifo_full       ),
        .empty              (wdata_fifo_empty      ),
        .valid              (wdata_fifo_valid      ),
        .prog_full_thresh   (10'd1023-FIFO_HEADROOM),
        .prog_full          (wdata_fifo_prog_full  )
    );

    /* araddr fifo (okFP -> MIG) */
    araddr_fifo_36_128 araddr_fifo (
        .rst                (fifo_rst              ),    // active-high
        .wr_clk             (okClk                 ),
        .rd_clk             (mig_clk               ),
        .din                (araddr_fifo_din       ),
        .wr_en              (araddr_fifo_wr_en     ),
        .rd_en              (araddr_fifo_rd_en     ),
        .dout               (araddr_fifo_dout      ),
        .full               (araddr_fifo_full      ),
        .empty              (araddr_fifo_empty     ),
        .valid              (araddr_fifo_valid     ),
        .prog_full_thresh   (7'd127-FIFO_HEADROOM  ),
        .prog_full          (araddr_fifo_prog_full )
    );

    /* rdata fifo (okFP <- MIG) */
    rdata_fifo_w256_128_r32_1024 rdata_fifo (
        .rst                (fifo_rst              ),    // active-high
        .wr_clk             (mig_clk               ),
        .rd_clk             (okClk                 ),
        .din                (rdata_fifo_din        ),
        .wr_en              (rdata_fifo_wr_en      ),
        .rd_en              (rdata_fifo_rd_en      ),
        .dout               (rdata_fifo_dout       ),
        .full               (rdata_fifo_full       ),
        .empty              (rdata_fifo_empty      ),
        .valid              (rdata_fifo_valid      ),
        .prog_full_thresh   (7'd127-FIFO_HEADROOM  ),
        .prog_full          (rdata_fifo_prog_full  )
    );


    always @(posedge mig_clk or negedge rstn) begin
        if (~rstn) begin
            mig_abort <= 1'b0;
        end
        else begin
            mig_abort <= abort;
        end
    end

    assign awaddr_fifo_wr_en       = (cmd_buf == CMD_DRAM_WRITE);    // We assumed awaddr_fifo will never be full
    assign awaddr_fifo_din         = {addr, axi_axlen};
    assign awaddr_fifo_rd_en       = axi_awready && (!awaddr_fifo_empty);
    assign {axi_awaddr, axi_awlen} = awaddr_fifo_rd_en && awaddr_fifo_valid ? awaddr_fifo_dout : 'd0;
    assign axi_awvalid             = awaddr_fifo_rd_en && awaddr_fifo_valid;


    assign wdata_fifo_wr_en        = pipe_in_valid;
    assign wdata_fifo_din          = pipe_din;
    assign wdata_fifo_rd_en        = axi_wready && (!wdata_fifo_empty);
    assign axi_wdata_pre_ord       = wdata_fifo_rd_en && wdata_fifo_valid ? wdata_fifo_dout : 'd0;
    assign axi_wdata               = reorder_4byte_blk(axi_wdata_pre_ord);
    assign axi_wvalid              = wdata_fifo_rd_en && wdata_fifo_valid;
    assign pipe_in_ready           = (state == S_DRAM_WRITE) && (!wdata_fifo_prog_full);


    assign araddr_fifo_wr_en       = (cmd_buf == CMD_DRAM_READ);    // We assumed araddr_fifo will never be full
    assign araddr_fifo_din         = {addr, axi_axlen};
    assign araddr_fifo_rd_en       = axi_arready && (!araddr_fifo_empty);
    assign {axi_araddr, axi_arlen} = araddr_fifo_rd_en && araddr_fifo_valid ? araddr_fifo_dout : 'd0;
    assign axi_arvalid             = araddr_fifo_rd_en && araddr_fifo_valid;


    assign rdata_fifo_wr_en        = axi_rvalid;
    assign axi_rdata_aft_ord       = reorder_4byte_blk(axi_rdata);
    assign rdata_fifo_din          = axi_rdata_aft_ord;

    assign rdata_fifo_rd_en        = (state == S_DRAM_READ) && (!rdata_fifo_empty) && pipe_out_ready_buf;
    assign pipe_dout               = rdata_fifo_valid ? rdata_fifo_dout : 'd0;
    assign pipe_out_valid          = rdata_fifo_valid;
    assign axi_rready              = !rdata_fifo_prog_full;



    //************************************************************
    // Instantiate FIFOs between okFP <-> Chip
    //************************************************************

    /* okFP -> Chip (start_net, single-rate, n_layers) */
    ok2chip_builtin_fifo_8_512 ok2chip_fifo (
        .rst                (fifo_rst              ),    // active-high
        .wr_clk             (okClk                 ),
        .rd_clk             (chip_clk              ),
        .din                (ok2chip_fifo_din      ),
        .wr_en              (ok2chip_fifo_wr_en    ),
        .rd_en              (ok2chip_fifo_rd_en    ),
        .dout               (ok2chip_fifo_dout     ),
        .full               (                      ),
        .empty              (ok2chip_fifo_empty    ),
        .valid              (ok2chip_fifo_valid    ),
        // .prog_full_thresh   (7'd127-FIFO_HEADROOM  ),
        .prog_full          (ok2chip_fifo_prog_full)
    );

    /* Chip -> okFP (done, clk_cnt) */
    chip2ok_builtin_fifo_32_512 chip2ok_fifo (
        .rst                (fifo_rst              ),    // active-high
        .wr_clk             (chip_clk              ),
        .rd_clk             (okClk                 ),
        .din                (chip2ok_fifo_din      ),
        .wr_en              (chip2ok_fifo_wr_en    ),
        .rd_en              (chip2ok_fifo_rd_en    ),
        .dout               (chip2ok_fifo_dout     ),
        .full               (                      ),
        .empty              (chip2ok_fifo_empty    ),
        .valid              (chip2ok_fifo_valid    ),
        // .prog_full_thresh   (7'd127-FIFO_HEADROOM  ),
        .prog_full          (chip2ok_fifo_prog_full)
    );

    assign ok2chip_fifo_wr_en = (cmd_buf == CMD_EXECUTE_NET);
    assign ok2chip_fifo_din   = {network_start, infinite_loop, n_layers};
    assign ok2chip_fifo_rd_en = ok2chip_fifo_valid;
    assign {chip_network_start, chip_infinite_loop, chip_n_layers} = ok2chip_fifo_valid ? ok2chip_fifo_dout : 8'd0;
    assign chip_single_rate = 1'b1;   // always 1'b1

    assign chip2ok_fifo_wr_en = chip_network_done;
    assign chip2ok_fifo_din   = {chip_network_done, chip_clk_cnt};
    assign chip2ok_fifo_rd_en = chip2ok_fifo_valid;
    assign {network_done, clk_cnt} = chip2ok_fifo_valid ? chip2ok_fifo_dout : 'd0;

    always @(posedge okClk) begin
        pipe_out_ready_buf <= pipe_out_ready;
    end

    reg [7:0] debug_chip_network_start_cnt;
    reg [7:0] debug_ok_network_start_cnt;
    reg [7:0] debug_chip_network_done_cnt;
    reg [7:0] debug_ok_network_done_cnt;

    assign ep39wire = {debug_chip_network_start_cnt, debug_ok_network_start_cnt, debug_chip_network_done_cnt, debug_ok_network_done_cnt};

    always @(posedge chip_clk or negedge rstn) begin
        if (~rstn) debug_chip_network_start_cnt <= 'd0;
        else if (chip_network_start) debug_chip_network_start_cnt <= debug_chip_network_start_cnt + 1;
    end

    always @(posedge okClk or negedge rstn) begin
        if (~rstn) debug_ok_network_start_cnt <= 'd0;
        else if (network_start) debug_ok_network_start_cnt <= debug_ok_network_start_cnt + 1;
    end

    always @(posedge chip_clk or negedge rstn) begin
        if (~rstn) debug_chip_network_done_cnt <= 'd0;
        else if (chip_network_done) debug_chip_network_done_cnt <= debug_chip_network_done_cnt + 1;
    end

    always @(posedge okClk or negedge rstn) begin
        if (~rstn) debug_ok_network_done_cnt <= 'd0;
        // else if (network_done) debug_ok_network_done_cnt <= debug_ok_network_done_cnt + 1;
        else if (network_done_buf) debug_ok_network_done_cnt <= debug_ok_network_done_cnt + 1;
    end



    //************************************************************
    // Signals for Debugging
    //************************************************************

    /* Debug */
    wire read_or_write;                // 0 for read, 1 for write
    wire [5:0] hist_idx;
    reg  [9:0] chip_clk_toggle_cnt;     // chip_clk domain
    reg  [9:0] chip_clk_toggle_cnt_ok;  // okClk domain

    reg  [3:0] ttf_axvalid_ok;

    assign read_or_write = ep05wire[0];
    assign hist_idx = ep06wire[5:0];
    // assign ep22wire = {done_cnt, start_cnt, arready_cnt, awready_cnt};


    assign ep24wire = read_or_write ? awaddr_hist[hist_idx] : araddr_hist[hist_idx];
    assign ep25wire = read_or_write ? awlen_hist[hist_idx] : arlen_hist[hist_idx];

    // assign {ep26wire, ep27wire, ep28wire, ep29wire, ep30wire, ep31wire, ep32wire, ep33wire} = rdata_hist[hist_idx];
    assign ep26wire = arvalid_cnt;
    assign ep27wire = rvalid_cnt;
    assign ep28wire = awvalid_cnt;
    assign ep29wire = wvalid_cnt;


    always @(posedge okClk or negedge rstn) begin
        if (~rstn) begin
            chip_clk_toggle_cnt_ok <= 'd0;
            ttf_axvalid_ok <= 'd0;
        end
        else begin
            chip_clk_toggle_cnt_ok <= chip_clk_toggle_cnt;
            ttf_axvalid_ok <= ttf_axvalid;
        end
    end

    always @(posedge chip_clk or negedge rstn) begin
        if (~rstn) begin
            chip_clk_toggle_cnt <= 'd0;
        end
        else begin
            if (chip_clk_toggle_cnt < 10'd1023)
                chip_clk_toggle_cnt <= chip_clk_toggle_cnt + 1;
        end
    end


    assign ep30wire = mig_rstate_cnt;
    assign ep31wire = mig_rvalid_cnt;
    assign ep32wire = mig_wstate_cnt;
    assign ep33wire = mig_wvalid_cnt;
    assign ep34wire = {28'd0, s_axi_wstate_debug, s_axi_wready_debug, s_axi_arready_debug, s_axi_rvalid_debug};
    // assign ep35wire = {mig_wstate_cnt, mig_rstate_cnt};
    assign ep36wire = {8'd0,
                       araddr_fifo_rd_en_debug, araddr_fifo_wr_en_debug, araddr_fifo_valid_debug, araddr_fifo_empty_debug, araddr_fifo_full_debug, araddr_fifo_prog_full_debug,
                       awaddr_fifo_rd_en_debug, awaddr_fifo_wr_en_debug, awaddr_fifo_valid_debug, awaddr_fifo_empty_debug, awaddr_fifo_full_debug, awaddr_fifo_prog_full_debug, 
                       rdata_fifo_rd_en_debug, rdata_fifo_wr_en_debug, rdata_fifo_valid_debug, rdata_fifo_empty_debug, rdata_fifo_full_debug, rdata_fifo_prog_full_debug, 
                       wdata_fifo_rd_en_debug, wdata_fifo_wr_en_debug, wdata_fifo_valid_debug, wdata_fifo_empty_debug, wdata_fifo_full_debug, wdata_fifo_prog_full_debug};

    assign ep37wire = ttf_axvalid_ok;

endmodule 


function [255:0] reorder_4byte_blk (
    input [255:0] data
);
    begin
        integer i;
        for (i = 0; i < 8; i = i + 1) begin
            reorder_4byte_blk[i*32 +: 32] = data[255 - i*32 -: 32];
        end
    end
endfunction